

module	GroundBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,	// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle,  //input that the pixel is within a bracket 

					output	logic	groundDR, 		//output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout   //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 


logic [0:14] [0:19]  MazeBiMapMask= 
{20'b	11111111111111111111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	11111111110000000001,
20'b	10000000000000001111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	10001111100000000001,
20'b	10000000000000000111,
20'b	10000000000000000001,
20'b	10000000000000000001,
20'b	11111111111111111111,
20'b	11111111111111111111};
 
 logic [0:1] [0:31] [0:31] [7:0]  object_colors  = {
{ {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h88,8'h40,8'h00,8'h00,8'h88,8'h00,8'h00,8'h80,8'h40,8'h00,8'h00,8'h80,8'h88,8'h00,8'h80,8'h80,8'h88,8'h00,8'h00,8'h40,8'h00,8'h40,8'h80,8'h80,8'h80,8'h88,8'h48,8'h10,8'h10,8'h00,8'h40},
	{8'h40,8'hc8,8'h40,8'h00,8'h00,8'h88,8'h40,8'h00,8'h80,8'h88,8'h00,8'h00,8'hc0,8'hc8,8'h00,8'h48,8'h88,8'h88,8'h40,8'h40,8'h40,8'h00,8'h48,8'h88,8'h88,8'hc0,8'hc0,8'h88,8'h10,8'h10,8'h00,8'h88},
	{8'h88,8'h88,8'h48,8'h10,8'h10,8'h48,8'hc8,8'h88,8'hc8,8'h88,8'h10,8'h10,8'hc8,8'h88,8'h50,8'h10,8'h08,8'h48,8'hc8,8'h88,8'h88,8'h50,8'h10,8'h08,8'h88,8'hc8,8'hc8,8'h88,8'h10,8'h18,8'h10,8'h88},
	{8'h50,8'h50,8'h10,8'h10,8'h10,8'h10,8'h50,8'h50,8'h50,8'h10,8'h10,8'h10,8'h50,8'h50,8'h10,8'h10,8'h10,8'h10,8'h50,8'h50,8'h50,8'h10,8'h10,8'h10,8'h10,8'h50,8'h50,8'h10,8'h10,8'h18,8'h10,8'h50},
	{8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h18,8'h10},
	{8'h10,8'h10,8'h10,8'h10,8'h10,8'h50,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h48,8'h48,8'h50,8'h10,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10},
	{8'h18,8'h10,8'h10,8'h10,8'h08,8'h88,8'h50,8'h10,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h88,8'hc8,8'h88,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10},
	{8'h10,8'h10,8'h18,8'h10,8'h10,8'h50,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18},
	{8'h10,8'h18,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h50,8'h50,8'h50,8'h50,8'h18,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h50,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h50},
	{8'h08,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h48,8'h88,8'h88,8'h48,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h48,8'h88,8'h50,8'h10,8'h10,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h88},
	{8'h50,8'h10,8'h18,8'h18,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h88},
	{8'h50,8'h10,8'h10,8'h18,8'h10,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h41},
	{8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h50,8'h50,8'h50,8'h10,8'h18,8'h18,8'h09},
	{8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h50,8'hc8,8'hc8,8'h88,8'h10,8'h18,8'h18,8'h10},
	{8'h10,8'h10,8'h10,8'h10,8'h10,8'h50,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h18,8'h10,8'h50,8'h50,8'h50,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h10,8'h10,8'h50,8'h10,8'h18,8'h18,8'h10,8'h88},
	{8'h50,8'h10,8'h10,8'h10,8'h08,8'h88,8'h50,8'h10,8'h18,8'h18,8'h18,8'h10,8'h10,8'h18,8'h10,8'h88,8'hc8,8'h88,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'hc8},
	{8'h50,8'h18,8'h10,8'h10,8'h10,8'h50,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'h10,8'h08,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h88,8'h88,8'h88,8'h50,8'h88},
	{8'h50,8'h10,8'h18,8'h10,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h48,8'h88,8'h50,8'h50,8'h48},
	{8'h50,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h50,8'h48,8'h48,8'h50,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h50,8'h50,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h09},
	{8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h08,8'h48,8'h50,8'h50,8'h18,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h50,8'h10,8'h18,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h88},
	{8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10,8'h18,8'h10,8'h18,8'h18,8'h18,8'h10,8'h10,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'h88},
	{8'h50,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h10,8'h18,8'h18,8'h18,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h50,8'hc8},
	{8'h50,8'h18,8'h18,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h48,8'h88,8'hc8,8'h10,8'h10,8'h18,8'h18,8'h10,8'h18,8'h18,8'h18,8'h50,8'h88,8'hc8,8'hc8,8'h50,8'h10,8'h48,8'hc8,8'hc8,8'h88,8'h50,8'hc8},
	{8'h50,8'h18,8'h10,8'h10,8'h10,8'h50,8'h10,8'h10,8'h10,8'h50,8'h88,8'h88,8'h10,8'h10,8'h10,8'h50,8'h50,8'h50,8'h10,8'h18,8'h10,8'h88,8'h88,8'h88,8'h50,8'h10,8'h10,8'h88,8'h88,8'h88,8'h50,8'h88},
	{8'h50,8'h10,8'h10,8'h10,8'h08,8'h88,8'h50,8'h18,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h10,8'h88,8'h88,8'h88,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h09},
	{8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h10,8'h18,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18},
	{8'h10,8'h10,8'h18,8'h18,8'h18,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h10,8'h10,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h10,8'h10,8'h10,8'h10,8'h10,8'h18,8'h18,8'h18,8'h18,8'h10,8'h48},
	{8'h88,8'h88,8'h50,8'h18,8'h10,8'h50,8'h88,8'h88,8'h88,8'h50,8'h10,8'h10,8'h90,8'h50,8'h10,8'h10,8'h10,8'h50,8'h88,8'h88,8'h50,8'h10,8'h10,8'h10,8'h50,8'h88,8'h88,8'h50,8'h10,8'h18,8'h10,8'hc8},
	{8'hc8,8'hc8,8'h88,8'h10,8'h50,8'h88,8'hc0,8'hc8,8'hc8,8'h88,8'h50,8'h50,8'hc8,8'hc8,8'h50,8'h10,8'h08,8'h48,8'hc8,8'hc8,8'h88,8'h50,8'h10,8'h08,8'h88,8'hc0,8'hc0,8'h88,8'h10,8'h10,8'h08,8'h88},
	{8'h01,8'h89,8'h41,8'h0a,8'h01,8'h89,8'h41,8'h02,8'h81,8'h89,8'h01,8'h41,8'h88,8'h89,8'h41,8'h89,8'h88,8'h89,8'h01,8'h01,8'h42,8'h01,8'h49,8'h88,8'h88,8'hc0,8'h88,8'h88,8'h10,8'h11,8'h09,8'h01},
	{8'h50,8'h18,8'h10,8'h10,8'h10,8'h50,8'h10,8'h10,8'h10,8'h50,8'h88,8'h88,8'h10,8'h10,8'h10,8'h50,8'h50,8'h50,8'h10,8'h18,8'h10,8'h88,8'h88,8'h88,8'h50,8'h10,8'h10,8'h88,8'h88,8'h88,8'h50,8'h88}
},
{	{8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h1b,8'h09,8'h09,8'h12},
	{8'h13,8'h12,8'h12,8'h12,8'h12,8'h0a,8'h09,8'h09,8'h09,8'h12,8'h12,8'h13,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h08,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h13,8'h0a,8'h12,8'h13},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h12,8'h12,8'h12,8'h13,8'h13,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h13,8'h13,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h0a,8'h13,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h11,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h08,8'h12,8'h12,8'h09},
	{8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h11,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h08,8'h12,8'h12,8'h09},
	{8'h09,8'h13,8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h13,8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h09,8'h09,8'h09,8'h09,8'h08,8'h12,8'h13,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h12,8'h0a,8'h0a,8'h12,8'h12,8'h13,8'h13,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h13,8'h0a,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h13,8'h0a,8'h09,8'h11,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h0a,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h09,8'h12,8'h09,8'h0a,8'h1b},
	{8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12},
	{8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h11,8'h12,8'h12,8'h09,8'h09,8'h09,8'h12,8'h12,8'h0a,8'h12,8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h12},
	{8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h13,8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12},
	{8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h13,8'h12,8'h09,8'h09,8'h09,8'h09,8'h13,8'h1b,8'h12,8'h13,8'h09,8'h09,8'h1b,8'h13,8'h13,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12},
	{8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h0a,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12},
	{8'h09,8'h09,8'h09,8'h13,8'h13,8'h13,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12},
	{8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h09,8'h09,8'h09},
	{8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h12,8'h12,8'h1b,8'h09,8'h09,8'h12},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h12,8'h12,8'h1b,8'h09,8'h09,8'h12},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h13,8'h12,8'h13,8'h12,8'h12,8'h0a,8'h12,8'h13,8'h13,8'h12,8'h12,8'h09,8'h08,8'h1b,8'h13,8'h13,8'h13,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h1b,8'h13,8'h09},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h11,8'h09,8'h11,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h13,8'h13,8'h0a},
	{8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h0a,8'h0a,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h0a,8'h12,8'h12,8'h12,8'h13,8'h13,8'h09},
	{8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h13,8'h13,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h12,8'h0a,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h13,8'h12,8'h09,8'h09,8'h12,8'h12,8'h13,8'h13,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h09},
	{8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h13,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h13},
	{8'h09,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h13,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h13,8'h13},
	{8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12},
	{8'h09,8'h12,8'h12,8'h09,8'h0a,8'h09,8'h09,8'h0a,8'h0a,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12},
	{8'h12,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h13,8'h12,8'h09,8'h09,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12},
	{8'h12,8'h09,8'h09,8'h09,8'h09,8'h13,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h0a,8'h09,8'h09,8'h12,8'h12,8'h12,8'h1a,8'h09,8'h0a,8'h12,8'h12,8'h09,8'h09,8'h09,8'h09,8'h09,8'h12,8'h12,8'h12}
 }
};

 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if ((InsideRectangle == 1'b1 )		& 								// only if inside the external bracket 
		   (MazeBiMapMask[offsetY[9:5] ][offsetX[9:5]] == 1'b1 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze 
				if(offsetY[8:5] == 0 || offsetY[8:5] == 14 || offsetX[9:5] == 0 || offsetX[9:5] == 19)
						RGBout <= object_colors[1][offsetY][offsetX] ;
				else
						RGBout <= object_colors[0][offsetY][offsetX] ;

		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign groundDR = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

